library verilog;
use verilog.vl_types.all;
entity Neural_network_TB is
end Neural_network_TB;
