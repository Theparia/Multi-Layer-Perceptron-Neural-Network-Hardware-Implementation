library verilog;
use verilog.vl_types.all;
entity Test_data_split is
    port(
        test_index      : in     vl_logic_vector(9 downto 0);
        \out\           : out    vl_logic_vector(495 downto 0)
    );
end Test_data_split;
